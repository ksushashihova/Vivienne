<svg width="144" height="45" viewBox="0 0 144 45" fill="none" xmlns="http://www.w3.org/2000/svg">
<path d="M11.0048 28.4286C14.5501 28.4286 17.4242 25.5545 17.4242 22.0092C17.4242 18.4639 14.5501 15.5899 11.0048 15.5899C7.45949 15.5899 4.58545 18.4639 4.58545 22.0092C4.58545 25.5545 7.45949 28.4286 11.0048 28.4286Z" fill="#F6D250"/>
<path d="M11.0045 32.0601C10.5002 32.0601 10.0875 31.6841 10.0875 31.1797V31.1064C10.0875 30.602 10.5002 30.1893 11.0045 30.1893C11.5089 30.1893 11.9216 30.602 11.9216 31.1064C11.9216 31.6107 11.5089 32.0601 11.0045 32.0601ZM17.5523 29.474C17.3139 29.474 17.0846 29.3823 16.9012 29.2081L16.782 29.0888C16.4243 28.7312 16.4243 28.1535 16.782 27.7958C17.1396 27.4382 17.7174 27.4382 18.075 27.7958L18.1942 27.915C18.5519 28.2727 18.5519 28.8504 18.1942 29.2081C18.02 29.3823 17.7907 29.474 17.5523 29.474ZM4.45681 29.474C4.21837 29.474 3.98911 29.3823 3.8057 29.2081C3.44805 28.8504 3.44805 28.2727 3.8057 27.915L3.92492 27.7958C4.28257 27.4382 4.86031 27.4382 5.21796 27.7958C5.57561 28.1535 5.57561 28.7312 5.21796 29.0888L5.09874 29.2081C4.9245 29.3823 4.68607 29.474 4.45681 29.474ZM20.1751 22.9263H20.1017C19.5973 22.9263 19.1846 22.5136 19.1846 22.0092C19.1846 21.5048 19.5973 21.0922 20.1017 21.0922C20.6061 21.0922 21.0554 21.5048 21.0554 22.0092C21.0554 22.5136 20.6794 22.9263 20.1751 22.9263ZM1.90741 22.9263H1.83404C1.32966 22.9263 0.916992 22.5136 0.916992 22.0092C0.916992 21.5048 1.32966 21.0922 1.83404 21.0922C2.33842 21.0922 2.78778 21.5048 2.78778 22.0092C2.78778 22.5136 2.41178 22.9263 1.90741 22.9263ZM17.4331 16.4977C17.1946 16.4977 16.9654 16.406 16.782 16.2318C16.4243 15.8741 16.4243 15.2964 16.782 14.9388L16.9012 14.8195C17.2588 14.4619 17.8366 14.4619 18.1942 14.8195C18.5519 15.1772 18.5519 15.7549 18.1942 16.1126L18.075 16.2318C17.9008 16.406 17.6715 16.4977 17.4331 16.4977ZM4.57602 16.4977C4.33759 16.4977 4.10833 16.406 3.92492 16.2318L3.8057 16.1034C3.44805 15.7458 3.44805 15.168 3.8057 14.8104C4.16335 14.4527 4.74109 14.4527 5.09874 14.8104L5.21796 14.9296C5.57561 15.2872 5.57561 15.865 5.21796 16.2226C5.04372 16.406 4.80529 16.4977 4.57602 16.4977ZM11.0045 13.7924C10.5002 13.7924 10.0875 13.4165 10.0875 12.9121V12.8387C10.0875 12.3343 10.5002 11.9217 11.0045 11.9217C11.5089 11.9217 11.9216 12.3343 11.9216 12.8387C11.9216 13.3431 11.5089 13.7924 11.0045 13.7924Z" fill="#F6D250"/>
<rect x="33.0137" width="77.0322" height="44.0184" rx="22.0092" fill="white"/>
<path d="M140.795 25.6132C140.648 25.3656 140.236 24.9804 139.208 25.1639C138.64 25.2647 138.062 25.3106 137.484 25.2831C135.348 25.1914 133.413 24.2101 132.065 22.697C130.872 21.3673 130.139 19.634 130.13 17.7633C130.13 16.7178 130.331 15.7091 130.744 14.7553C131.148 13.8291 130.863 13.3431 130.662 13.1413C130.451 12.9304 129.955 12.6369 128.983 13.0405C125.233 14.6178 122.912 18.3777 123.188 22.4035C123.463 26.191 126.122 29.4281 129.644 30.6478C130.487 30.9413 131.377 31.1155 132.294 31.1522C132.441 31.1614 132.587 31.1705 132.734 31.1705C135.806 31.1705 138.686 29.7216 140.501 27.2547C141.116 26.4019 140.951 25.8608 140.795 25.6132Z" fill="#0088FF"/>
</svg>
